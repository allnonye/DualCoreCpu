`timescale 1ns / 1ps


module SevsegDisplay(
      input [3:0] Dig0,
      input [3:0] Dig1,
      input [3:0] Dig2,
      input [3:0] Dig3,
      input Cin,
      input clr,
      input clk,
      output [3:0] AN,
      output [6:0] CA
    );
    
  //  Sevseg s0 (.DigA(Dig0), .DigB(Dig1), .DigC(Dig2), .DigD(Dig3), .Cin(Cin), .clr(clr), .clk(clk), .AN(AN), .CA(C
    
    
endmodule
